*XOR Gate using Transmission gate:
.include "D:\mosmodel.txt"
 VDD 1 0 1.8V
 Va 2 0 PULSE 0 1.8 0 1n 1n 10u 20u
 Vb 4 0 PULSE 0 1.8 0 1n 1n 20u 40u
 Cl 6 0 100f
.model mn NMOS L=0.18u W=0.36u
.model mp PMOS L=0.18u W=0.72u
 M1 3 2 1 1 mp AS = 0.648p AD = 0.648p PS = 3.24u PD = 3.24u
 M2 3 2 0 0 mn AS = 0.648p AD = 0.648p PS = 3.24u PD = 3.24u
 M3 5 4 1 1 mp AS = 0.648p AD = 0.648p PS = 3.24u PD = 3.24u
 M4 5 4 0 0 mn AS = 0.648p AD = 0.648p PS = 3.24u PD = 3.24u
 M5 6 2 4 1 mp AS = 0.648p AD = 0.648p PS = 3.24u PD = 3.24u
 M6 6 3 4 0 mn AS = 0.648p AD = 0.648p PS = 3.24u PD = 3.24u
 M7 6 3 5 1 mp AS = 0.648p AD = 0.648p PS = 3.24u PD = 3.24u
 M8 6 2 5 0 mn AS = 0.648p AD = 0.648p PS = 3.24u PD = 3.24u
.TRAN 1u 80u
.PROBE
.END
